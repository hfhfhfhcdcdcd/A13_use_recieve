module  use_recieve(
    input rst,
    input sclk,
    input [7:0]data,
    input rx_done,
    output [7:0]ctrl,
    output [31:0]time_ctrl
);
/*
�ƶ�һ��Э�飺�����������֣���������ģ��������У�
��һ������������һģ�� ctrl �˿ڵġ���Щ��������
����һģ��� time_ctrl �˿ڵġ�

Լ���������յ�rx_done�ź�ʱ����ʼ��⴫����������ݡ�
����Э������ǣ�����⵽rx_done�ź�ʱ���ȿ����Ƿ�
���������ݣ�oxAB��oxCD, �����⵽���������ݣ���ʼ
���մ����������ݡ����Ʋ���40bit����Ϊ��һ��ģ��Ҫ�õ�
40bit��8bitctrl��32bittime_ctrl���������꣬�����Ȼ
Ҫ����Ƿ���oxEF����ֽڣ��еĻ�˵���ղŽ��յ�������
����ȷ�ģ�û�������øղŽ��յ������ݡ�

��ȻҪ
*/

endmodule